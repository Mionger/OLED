module SPI
(
    
);

endmodule