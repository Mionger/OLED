module  Divider
(
    DI,
    DO,
    N
);
    input DI;
    input N;

    output DO;

    reg DO = 0;

    integer t_cnt = 0;
    always @(posedge DI) begin
        if(t_cnt<N/2-1) begin
            t_cnt <= t_cnt + 1;
        end
        else begin
            t_cnt <= 0;
            DO    <= ~DO;
        end
    end
endmodule